package wrapper_shared_pkg;
int error_count;
int correct_count;
int error_count_2;
int correct_count_2;
int error_count_r;
int correct_count_r;
int error_count_w;
int correct_count_w;
int error_count_s;
int correct_count_s;
int error_count_2_s;
int correct_count_2_s;
int Count_seq, i, address_recieved;
int count;
bit start_read;

endpackage